module check

struct Settings {
}
