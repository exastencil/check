module check

pub struct Settings {
	store_path string
}
