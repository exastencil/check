module check

pub struct Settings {
pub:
	store_path string
}
