module web

struct Feed {
	url string
}
