module twitter

struct Account {
	handle   string
	password string
}
