module mail

struct Account {
	address  string
	password string
	imap     string
}
